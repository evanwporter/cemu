`ifndef PPU_TYPES_SV
`define PPU_TYPES_SV 

typedef enum logic [1:0] {
  PPU_MODE_0,
  PPU_MODE_1,
  PPU_MODE_2,
  PPU_MODE_3
} ppu_mode_t;

`endif  // PPU_TYPES_SV
