package gb_types_pkg;

  typedef enum logic [1:0] {
    T1,
    T2,
    T3,
    T4
  } t_phase_t;

endpackage : gb_types_pkg
