`ifndef MMU_TYPES_SV
`define MMU_TYPES_SV 

typedef logic [15:0] address_t;

`endif
