package gba_types_pkg;
  typedef logic [31:0] word_t;

  typedef logic [15:0] half_t;

  typedef logic [7:0] byte_t;

endpackage : gba_types_pkg
