`include "ppu/fetcher/Fetcher.sv"
`include "ppu/fifo/FIFO.sv"
`include "ppu/Framebuffer.sv"
`include "ppu/fetcher/ObjFetcher.sv"
`include "ppu/fifo/ObjFIFO.sv"
`include "ppu/PPU.sv"

import ppu_types_pkg::*;
import ppu_util_pkg::*;

module ppu_top (
    input logic clk,
    input logic reset
);

  GB_Bus_if ppu_bus ();
  GB_Interrupt_if IF_bus ();
  GB_DMA_if dma_bus ();

  GB_PPU ppu (
      clk,
      reset,
      ppu_bus,
      IF_bus,
      dma_bus
  );

  initial begin
    ppu.regs.SCX  = 8'd0;
    ppu.regs.SCY  = 8'd0;
    ppu.regs.LCDC = 8'b1001_0001;  // LCD on, BG on, 0x8000 tiles, 0x9800 map

    ppu.VRAM <= '{default: 8'h00};

    ppu.mode = PPU_MODE_3;
  end

endmodule
