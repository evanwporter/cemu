package ppu_fetcher_types_pkg;

  typedef enum logic {
    DOT_PHASE_0,
    DOT_PHASE_1
  } dot_phase_t;

endpackage : ppu_fetcher_types_pkg

