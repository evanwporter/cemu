module ALU (
    input logic clk,
    input logic reset
);


endmodule : ALU
