// From the Gearboy emulator
localparam logic [7:0] BOOT_DMG[0:255] = '{
    8'h31,
    8'hFE,
    8'hFF,
    8'hAF,
    8'h21,
    8'hFF,
    8'h9F,
    8'h32,
    8'hCB,
    8'h7C,
    8'h20,
    8'hFB,
    8'h21,
    8'h26,
    8'hFF,
    8'h0E,
    8'h11,
    8'h3E,
    8'h80,
    8'h32,
    8'hE2,
    8'h0C,
    8'h3E,
    8'hF3,
    8'hE2,
    8'h32,
    8'h3E,
    8'h77,
    8'h77,
    8'h3E,
    8'hFC,
    8'hE0,
    8'h47,
    8'h11,
    8'h04,
    8'h01,
    8'h21,
    8'h10,
    8'h80,
    8'h1A,
    8'hCD,
    8'h95,
    8'h00,
    8'hCD,
    8'h96,
    8'h00,
    8'h13,
    8'h7B,
    8'hFE,
    8'h34,
    8'h20,
    8'hF3,
    8'h11,
    8'hD8,
    8'h00,
    8'h06,
    8'h08,
    8'h1A,
    8'h13,
    8'h22,
    8'h23,
    8'h05,
    8'h20,
    8'hF9,
    8'h3E,
    8'h19,
    8'hEA,
    8'h10,
    8'h99,
    8'h21,
    8'h2F,
    8'h99,
    8'h0E,
    8'h0C,
    8'h3D,
    8'h28,
    8'h08,
    8'h32,
    8'h0D,
    8'h20,
    8'hF9,
    8'h2E,
    8'h0F,
    8'h18,
    8'hF3,
    8'h67,
    8'h3E,
    8'h64,
    8'h57,
    8'hE0,
    8'h42,
    8'h3E,
    8'h91,
    8'hE0,
    8'h40,
    8'h04,
    8'h1E,
    8'h02,
    8'h0E,
    8'h0C,
    8'hF0,
    8'h44,
    8'hFE,
    8'h90,
    8'h20,
    8'hFA,
    8'h0D,
    8'h20,
    8'hF7,
    8'h1D,
    8'h20,
    8'hF2,
    8'h0E,
    8'h13,
    8'h24,
    8'h7C,
    8'h1E,
    8'h83,
    8'hFE,
    8'h62,
    8'h28,
    8'h06,
    8'h1E,
    8'hC1,
    8'hFE,
    8'h64,
    8'h20,
    8'h06,
    8'h7B,
    8'hE2,
    8'h0C,
    8'h3E,
    8'h87,
    8'hE2,
    8'hF0,
    8'h42,
    8'h90,
    8'hE0,
    8'h42,
    8'h15,
    8'h20,
    8'hD2,
    8'h05,
    8'h20,
    8'h4F,
    8'h16,
    8'h20,
    8'h18,
    8'hCB,
    8'h4F,
    8'h06,
    8'h04,
    8'hC5,
    8'hCB,
    8'h11,
    8'h17,
    8'hC1,
    8'hCB,
    8'h11,
    8'h17,
    8'h05,
    8'h20,
    8'hF5,
    8'h22,
    8'h23,
    8'h22,
    8'h23,
    8'hC9,
    8'hCE,
    8'hED,
    8'h66,
    8'h66,
    8'hCC,
    8'h0D,
    8'h00,
    8'h0B,
    8'h03,
    8'h73,
    8'h00,
    8'h83,
    8'h00,
    8'h0C,
    8'h00,
    8'h0D,
    8'h00,
    8'h08,
    8'h11,
    8'h1F,
    8'h88,
    8'h89,
    8'h00,
    8'h0E,
    8'hDC,
    8'hCC,
    8'h6E,
    8'hE6,
    8'hDD,
    8'hDD,
    8'hD9,
    8'h99,
    8'hBB,
    8'hBB,
    8'h67,
    8'h63,
    8'h6E,
    8'h0E,
    8'hEC,
    8'hCC,
    8'hDD,
    8'hDC,
    8'h99,
    8'h9F,
    8'hBB,
    8'hB9,
    8'h33,
    8'h3E,
    8'h3C,
    8'h42,
    8'hB9,
    8'hA5,
    8'hB9,
    8'hA5,
    8'h42,
    8'h3C,
    8'h21,
    8'h04,
    8'h01,
    8'h11,
    8'hA8,
    8'h00,
    8'h1A,
    8'h13,
    8'hBE,
    8'h00,
    8'h00,
    8'h23,
    8'h7D,
    8'hFE,
    8'h34,
    8'h20,
    8'hF5,
    8'h06,
    8'h19,
    8'h78,
    8'h86,
    8'h23,
    8'h05,
    8'h20,
    8'hFB,
    8'h86,
    8'h00,
    8'h00,
    8'h3E,
    8'h01,
    8'hE0,
    8'h50
};
